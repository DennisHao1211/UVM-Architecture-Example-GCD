/nethome/hhao40/uvm_onboarding/src/uvm/tests/gcd_test_pkg.sv