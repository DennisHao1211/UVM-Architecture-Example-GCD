/nethome/hhao40/uvm_onboarding/src/uvm/agent/gcd_monitor.sv