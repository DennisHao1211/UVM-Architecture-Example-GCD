/nethome/hhao40/uvm_onboarding/src/uvm/env/gcd_sb.sv