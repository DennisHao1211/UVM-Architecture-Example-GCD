/nethome/hhao40/uvm_onboarding/src/uvm/env/gcd_env_pkg.sv