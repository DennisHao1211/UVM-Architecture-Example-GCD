/nethome/hhao40/uvm_onboarding/src/uvm/sequences/gcd_sequence.svh