/nethome/hhao40/uvm_onboarding/src/uvm/tests/gcd_base_test.svh