/nethome/hhao40/uvm_onboarding/src/sv/rtl/gcd_pkg.sv