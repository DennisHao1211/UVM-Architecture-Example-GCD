/nethome/hhao40/uvm_onboarding/src/uvm/tb/gcd_if.sv