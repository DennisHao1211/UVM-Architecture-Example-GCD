/nethome/hhao40/uvm_onboarding/src/uvm/sequences/gcd_seq_pkg.sv